module E(input [1:32] in, output [1:48] out);
  assign out[1] = in[32];
  assign out[2] = in[1];
  assign out[3] = in[2];
  assign out[4] = in[3];
  assign out[5] = in[4];
  assign out[6] = in[5];
  assign out[7] = in[4];
  assign out[8] = in[5];
  assign out[9] = in[6];
  assign out[10] = in[7];
  assign out[11] = in[8];
  assign out[12] = in[9];
  assign out[13] = in[8];
  assign out[14] = in[9];
  assign out[15] = in[10];
  assign out[16] = in[11];
  assign out[17] = in[12];
  assign out[18] = in[13];
  assign out[19] = in[12];
  assign out[20] = in[13];
  assign out[21] = in[14];
  assign out[22] = in[15];
  assign out[23] = in[16];
  assign out[24] = in[17];
  assign out[25] = in[16];
  assign out[26] = in[17];
  assign out[27] = in[18];
  assign out[28] = in[19];
  assign out[29] = in[20];
  assign out[30] = in[21];
  assign out[31] = in[20];
  assign out[32] = in[21];
  assign out[33] = in[22];
  assign out[34] = in[23];
  assign out[35] = in[24];
  assign out[36] = in[25];
  assign out[37] = in[24];
  assign out[38] = in[25];
  assign out[39] = in[26];
  assign out[40] = in[27];
  assign out[41] = in[28];
  assign out[42] = in[29];
  assign out[43] = in[28];
  assign out[44] = in[29];
  assign out[45] = in[30];
  assign out[46] = in[31];
  assign out[47] = in[32];
  assign out[48] = in[1];
endmodule
module P(input [1:32] in, output [1:32] out);
  assign out[1] = in[16];
  assign out[2] = in[7];
  assign out[3] = in[20];
  assign out[4] = in[21];
  assign out[5] = in[29];
  assign out[6] = in[12];
  assign out[7] = in[28];
  assign out[8] = in[17];
  assign out[9] = in[1];
  assign out[10] = in[15];
  assign out[11] = in[23];
  assign out[12] = in[26];
  assign out[13] = in[5];
  assign out[14] = in[18];
  assign out[15] = in[31];
  assign out[16] = in[10];
  assign out[17] = in[2];
  assign out[18] = in[8];
  assign out[19] = in[24];
  assign out[20] = in[14];
  assign out[21] = in[32];
  assign out[22] = in[27];
  assign out[23] = in[3];
  assign out[24] = in[9];
  assign out[25] = in[19];
  assign out[26] = in[13];
  assign out[27] = in[30];
  assign out[28] = in[6];
  assign out[29] = in[22];
  assign out[30] = in[11];
  assign out[31] = in[4];
  assign out[32] = in[25];
endmodule
module S1(input [6:1] in, output reg [4:1] out);
  always @* case (in)
    0 : out = 14;
    1 : out = 0;
    2 : out = 4;
    3 : out = 15;
    4 : out = 13;
    5 : out = 7;
    6 : out = 1;
    7 : out = 4;
    8 : out = 2;
    9 : out = 14;
    10 : out = 15;
    11 : out = 2;
    12 : out = 11;
    13 : out = 13;
    14 : out = 8;
    15 : out = 1;
    16 : out = 3;
    17 : out = 10;
    18 : out = 10;
    19 : out = 6;
    20 : out = 6;
    21 : out = 12;
    22 : out = 12;
    23 : out = 11;
    24 : out = 5;
    25 : out = 9;
    26 : out = 9;
    27 : out = 5;
    28 : out = 0;
    29 : out = 3;
    30 : out = 7;
    31 : out = 8;
    32 : out = 4;
    33 : out = 15;
    34 : out = 1;
    35 : out = 12;
    36 : out = 14;
    37 : out = 8;
    38 : out = 8;
    39 : out = 2;
    40 : out = 13;
    41 : out = 4;
    42 : out = 6;
    43 : out = 9;
    44 : out = 2;
    45 : out = 1;
    46 : out = 11;
    47 : out = 7;
    48 : out = 15;
    49 : out = 5;
    50 : out = 12;
    51 : out = 11;
    52 : out = 9;
    53 : out = 3;
    54 : out = 7;
    55 : out = 14;
    56 : out = 3;
    57 : out = 10;
    58 : out = 10;
    59 : out = 0;
    60 : out = 5;
    61 : out = 6;
    62 : out = 0;
    63 : out = 13;
  endcase
endmodule
module S2(input [6:1] in, output reg [4:1] out);
  always @* case (in)
    0 : out = 15;
    1 : out = 3;
    2 : out = 1;
    3 : out = 13;
    4 : out = 8;
    5 : out = 4;
    6 : out = 14;
    7 : out = 7;
    8 : out = 6;
    9 : out = 15;
    10 : out = 11;
    11 : out = 2;
    12 : out = 3;
    13 : out = 8;
    14 : out = 4;
    15 : out = 14;
    16 : out = 9;
    17 : out = 12;
    18 : out = 7;
    19 : out = 0;
    20 : out = 2;
    21 : out = 1;
    22 : out = 13;
    23 : out = 10;
    24 : out = 12;
    25 : out = 6;
    26 : out = 0;
    27 : out = 9;
    28 : out = 5;
    29 : out = 11;
    30 : out = 10;
    31 : out = 5;
    32 : out = 0;
    33 : out = 13;
    34 : out = 14;
    35 : out = 8;
    36 : out = 7;
    37 : out = 10;
    38 : out = 11;
    39 : out = 1;
    40 : out = 10;
    41 : out = 3;
    42 : out = 4;
    43 : out = 15;
    44 : out = 13;
    45 : out = 4;
    46 : out = 1;
    47 : out = 2;
    48 : out = 5;
    49 : out = 11;
    50 : out = 8;
    51 : out = 6;
    52 : out = 12;
    53 : out = 7;
    54 : out = 6;
    55 : out = 12;
    56 : out = 9;
    57 : out = 0;
    58 : out = 3;
    59 : out = 5;
    60 : out = 2;
    61 : out = 14;
    62 : out = 15;
    63 : out = 9;
  endcase
endmodule
module S3(input [6:1] in, output reg [4:1] out);
  always @* case (in)
    0 : out = 10;
    1 : out = 13;
    2 : out = 0;
    3 : out = 7;
    4 : out = 9;
    5 : out = 0;
    6 : out = 14;
    7 : out = 9;
    8 : out = 6;
    9 : out = 3;
    10 : out = 3;
    11 : out = 4;
    12 : out = 15;
    13 : out = 6;
    14 : out = 5;
    15 : out = 10;
    16 : out = 1;
    17 : out = 2;
    18 : out = 13;
    19 : out = 8;
    20 : out = 12;
    21 : out = 5;
    22 : out = 7;
    23 : out = 14;
    24 : out = 11;
    25 : out = 12;
    26 : out = 4;
    27 : out = 11;
    28 : out = 2;
    29 : out = 15;
    30 : out = 8;
    31 : out = 1;
    32 : out = 13;
    33 : out = 1;
    34 : out = 6;
    35 : out = 10;
    36 : out = 4;
    37 : out = 13;
    38 : out = 9;
    39 : out = 0;
    40 : out = 8;
    41 : out = 6;
    42 : out = 15;
    43 : out = 9;
    44 : out = 3;
    45 : out = 8;
    46 : out = 0;
    47 : out = 7;
    48 : out = 11;
    49 : out = 4;
    50 : out = 1;
    51 : out = 15;
    52 : out = 2;
    53 : out = 14;
    54 : out = 12;
    55 : out = 3;
    56 : out = 5;
    57 : out = 11;
    58 : out = 10;
    59 : out = 5;
    60 : out = 14;
    61 : out = 2;
    62 : out = 7;
    63 : out = 12;
  endcase
endmodule
module S4(input [6:1] in, output reg [4:1] out);
  always @* case (in)
    0 : out = 7;
    1 : out = 13;
    2 : out = 13;
    3 : out = 8;
    4 : out = 14;
    5 : out = 11;
    6 : out = 3;
    7 : out = 5;
    8 : out = 0;
    9 : out = 6;
    10 : out = 6;
    11 : out = 15;
    12 : out = 9;
    13 : out = 0;
    14 : out = 10;
    15 : out = 3;
    16 : out = 1;
    17 : out = 4;
    18 : out = 2;
    19 : out = 7;
    20 : out = 8;
    21 : out = 2;
    22 : out = 5;
    23 : out = 12;
    24 : out = 11;
    25 : out = 1;
    26 : out = 12;
    27 : out = 10;
    28 : out = 4;
    29 : out = 14;
    30 : out = 15;
    31 : out = 9;
    32 : out = 10;
    33 : out = 3;
    34 : out = 6;
    35 : out = 15;
    36 : out = 9;
    37 : out = 0;
    38 : out = 0;
    39 : out = 6;
    40 : out = 12;
    41 : out = 10;
    42 : out = 11;
    43 : out = 1;
    44 : out = 7;
    45 : out = 13;
    46 : out = 13;
    47 : out = 8;
    48 : out = 15;
    49 : out = 9;
    50 : out = 1;
    51 : out = 4;
    52 : out = 3;
    53 : out = 5;
    54 : out = 14;
    55 : out = 11;
    56 : out = 5;
    57 : out = 12;
    58 : out = 2;
    59 : out = 7;
    60 : out = 8;
    61 : out = 2;
    62 : out = 4;
    63 : out = 14;
  endcase
endmodule
module S5(input [6:1] in, output reg [4:1] out);
  always @* case (in)
    0 : out = 2;
    1 : out = 14;
    2 : out = 12;
    3 : out = 11;
    4 : out = 4;
    5 : out = 2;
    6 : out = 1;
    7 : out = 12;
    8 : out = 7;
    9 : out = 4;
    10 : out = 10;
    11 : out = 7;
    12 : out = 11;
    13 : out = 13;
    14 : out = 6;
    15 : out = 1;
    16 : out = 8;
    17 : out = 5;
    18 : out = 5;
    19 : out = 0;
    20 : out = 3;
    21 : out = 15;
    22 : out = 15;
    23 : out = 10;
    24 : out = 13;
    25 : out = 3;
    26 : out = 0;
    27 : out = 9;
    28 : out = 14;
    29 : out = 8;
    30 : out = 9;
    31 : out = 6;
    32 : out = 4;
    33 : out = 11;
    34 : out = 2;
    35 : out = 8;
    36 : out = 1;
    37 : out = 12;
    38 : out = 11;
    39 : out = 7;
    40 : out = 10;
    41 : out = 1;
    42 : out = 13;
    43 : out = 14;
    44 : out = 7;
    45 : out = 2;
    46 : out = 8;
    47 : out = 13;
    48 : out = 15;
    49 : out = 6;
    50 : out = 9;
    51 : out = 15;
    52 : out = 12;
    53 : out = 0;
    54 : out = 5;
    55 : out = 9;
    56 : out = 6;
    57 : out = 10;
    58 : out = 3;
    59 : out = 4;
    60 : out = 0;
    61 : out = 5;
    62 : out = 14;
    63 : out = 3;
  endcase
endmodule
module S6(input [6:1] in, output reg [4:1] out);
  always @* case (in)
    0 : out = 12;
    1 : out = 10;
    2 : out = 1;
    3 : out = 15;
    4 : out = 10;
    5 : out = 4;
    6 : out = 15;
    7 : out = 2;
    8 : out = 9;
    9 : out = 7;
    10 : out = 2;
    11 : out = 12;
    12 : out = 6;
    13 : out = 9;
    14 : out = 8;
    15 : out = 5;
    16 : out = 0;
    17 : out = 6;
    18 : out = 13;
    19 : out = 1;
    20 : out = 3;
    21 : out = 13;
    22 : out = 4;
    23 : out = 14;
    24 : out = 14;
    25 : out = 0;
    26 : out = 7;
    27 : out = 11;
    28 : out = 5;
    29 : out = 3;
    30 : out = 11;
    31 : out = 8;
    32 : out = 9;
    33 : out = 4;
    34 : out = 14;
    35 : out = 3;
    36 : out = 15;
    37 : out = 2;
    38 : out = 5;
    39 : out = 12;
    40 : out = 2;
    41 : out = 9;
    42 : out = 8;
    43 : out = 5;
    44 : out = 12;
    45 : out = 15;
    46 : out = 3;
    47 : out = 10;
    48 : out = 7;
    49 : out = 11;
    50 : out = 0;
    51 : out = 14;
    52 : out = 4;
    53 : out = 1;
    54 : out = 10;
    55 : out = 7;
    56 : out = 1;
    57 : out = 6;
    58 : out = 13;
    59 : out = 0;
    60 : out = 11;
    61 : out = 8;
    62 : out = 6;
    63 : out = 13;
  endcase
endmodule
module S7(input [6:1] in, output reg [4:1] out);
  always @* case (in)
    0 : out = 4;
    1 : out = 13;
    2 : out = 11;
    3 : out = 0;
    4 : out = 2;
    5 : out = 11;
    6 : out = 14;
    7 : out = 7;
    8 : out = 15;
    9 : out = 4;
    10 : out = 0;
    11 : out = 9;
    12 : out = 8;
    13 : out = 1;
    14 : out = 13;
    15 : out = 10;
    16 : out = 3;
    17 : out = 14;
    18 : out = 12;
    19 : out = 3;
    20 : out = 9;
    21 : out = 5;
    22 : out = 7;
    23 : out = 12;
    24 : out = 5;
    25 : out = 2;
    26 : out = 10;
    27 : out = 15;
    28 : out = 6;
    29 : out = 8;
    30 : out = 1;
    31 : out = 6;
    32 : out = 1;
    33 : out = 6;
    34 : out = 4;
    35 : out = 11;
    36 : out = 11;
    37 : out = 13;
    38 : out = 13;
    39 : out = 8;
    40 : out = 12;
    41 : out = 1;
    42 : out = 3;
    43 : out = 4;
    44 : out = 7;
    45 : out = 10;
    46 : out = 14;
    47 : out = 7;
    48 : out = 10;
    49 : out = 9;
    50 : out = 15;
    51 : out = 5;
    52 : out = 6;
    53 : out = 0;
    54 : out = 8;
    55 : out = 15;
    56 : out = 0;
    57 : out = 14;
    58 : out = 5;
    59 : out = 2;
    60 : out = 9;
    61 : out = 3;
    62 : out = 2;
    63 : out = 12;
  endcase
endmodule
module S8(input [6:1] in, output reg [4:1] out);
  always @* case (in)
    0 : out = 13;
    1 : out = 1;
    2 : out = 2;
    3 : out = 15;
    4 : out = 8;
    5 : out = 13;
    6 : out = 4;
    7 : out = 8;
    8 : out = 6;
    9 : out = 10;
    10 : out = 15;
    11 : out = 3;
    12 : out = 11;
    13 : out = 7;
    14 : out = 1;
    15 : out = 4;
    16 : out = 10;
    17 : out = 12;
    18 : out = 9;
    19 : out = 5;
    20 : out = 3;
    21 : out = 6;
    22 : out = 14;
    23 : out = 11;
    24 : out = 5;
    25 : out = 0;
    26 : out = 0;
    27 : out = 14;
    28 : out = 12;
    29 : out = 9;
    30 : out = 7;
    31 : out = 2;
    32 : out = 7;
    33 : out = 2;
    34 : out = 11;
    35 : out = 1;
    36 : out = 4;
    37 : out = 14;
    38 : out = 1;
    39 : out = 7;
    40 : out = 9;
    41 : out = 4;
    42 : out = 12;
    43 : out = 10;
    44 : out = 14;
    45 : out = 8;
    46 : out = 2;
    47 : out = 13;
    48 : out = 0;
    49 : out = 15;
    50 : out = 6;
    51 : out = 12;
    52 : out = 10;
    53 : out = 9;
    54 : out = 13;
    55 : out = 0;
    56 : out = 15;
    57 : out = 3;
    58 : out = 3;
    59 : out = 5;
    60 : out = 5;
    61 : out = 6;
    62 : out = 8;
    63 : out = 11;
  endcase
endmodule
module IP(input [1:64] in, output [1:64] out);
  assign out[1] = in[58];
  assign out[2] = in[50];
  assign out[3] = in[42];
  assign out[4] = in[34];
  assign out[5] = in[26];
  assign out[6] = in[18];
  assign out[7] = in[10];
  assign out[8] = in[2];
  assign out[9] = in[60];
  assign out[10] = in[52];
  assign out[11] = in[44];
  assign out[12] = in[36];
  assign out[13] = in[28];
  assign out[14] = in[20];
  assign out[15] = in[12];
  assign out[16] = in[4];
  assign out[17] = in[62];
  assign out[18] = in[54];
  assign out[19] = in[46];
  assign out[20] = in[38];
  assign out[21] = in[30];
  assign out[22] = in[22];
  assign out[23] = in[14];
  assign out[24] = in[6];
  assign out[25] = in[64];
  assign out[26] = in[56];
  assign out[27] = in[48];
  assign out[28] = in[40];
  assign out[29] = in[32];
  assign out[30] = in[24];
  assign out[31] = in[16];
  assign out[32] = in[8];
  assign out[33] = in[57];
  assign out[34] = in[49];
  assign out[35] = in[41];
  assign out[36] = in[33];
  assign out[37] = in[25];
  assign out[38] = in[17];
  assign out[39] = in[9];
  assign out[40] = in[1];
  assign out[41] = in[59];
  assign out[42] = in[51];
  assign out[43] = in[43];
  assign out[44] = in[35];
  assign out[45] = in[27];
  assign out[46] = in[19];
  assign out[47] = in[11];
  assign out[48] = in[3];
  assign out[49] = in[61];
  assign out[50] = in[53];
  assign out[51] = in[45];
  assign out[52] = in[37];
  assign out[53] = in[29];
  assign out[54] = in[21];
  assign out[55] = in[13];
  assign out[56] = in[5];
  assign out[57] = in[63];
  assign out[58] = in[55];
  assign out[59] = in[47];
  assign out[60] = in[39];
  assign out[61] = in[31];
  assign out[62] = in[23];
  assign out[63] = in[15];
  assign out[64] = in[7];
endmodule
module IP_inv(input [1:64] in, output [1:64] out);
  assign out[1] = in[40];
  assign out[2] = in[8];
  assign out[3] = in[48];
  assign out[4] = in[16];
  assign out[5] = in[56];
  assign out[6] = in[24];
  assign out[7] = in[64];
  assign out[8] = in[32];
  assign out[9] = in[39];
  assign out[10] = in[7];
  assign out[11] = in[47];
  assign out[12] = in[15];
  assign out[13] = in[55];
  assign out[14] = in[23];
  assign out[15] = in[63];
  assign out[16] = in[31];
  assign out[17] = in[38];
  assign out[18] = in[6];
  assign out[19] = in[46];
  assign out[20] = in[14];
  assign out[21] = in[54];
  assign out[22] = in[22];
  assign out[23] = in[62];
  assign out[24] = in[30];
  assign out[25] = in[37];
  assign out[26] = in[5];
  assign out[27] = in[45];
  assign out[28] = in[13];
  assign out[29] = in[53];
  assign out[30] = in[21];
  assign out[31] = in[61];
  assign out[32] = in[29];
  assign out[33] = in[36];
  assign out[34] = in[4];
  assign out[35] = in[44];
  assign out[36] = in[12];
  assign out[37] = in[52];
  assign out[38] = in[20];
  assign out[39] = in[60];
  assign out[40] = in[28];
  assign out[41] = in[35];
  assign out[42] = in[3];
  assign out[43] = in[43];
  assign out[44] = in[11];
  assign out[45] = in[51];
  assign out[46] = in[19];
  assign out[47] = in[59];
  assign out[48] = in[27];
  assign out[49] = in[34];
  assign out[50] = in[2];
  assign out[51] = in[42];
  assign out[52] = in[10];
  assign out[53] = in[50];
  assign out[54] = in[18];
  assign out[55] = in[58];
  assign out[56] = in[26];
  assign out[57] = in[33];
  assign out[58] = in[1];
  assign out[59] = in[41];
  assign out[60] = in[9];
  assign out[61] = in[49];
  assign out[62] = in[17];
  assign out[63] = in[57];
  assign out[64] = in[25];
endmodule
module PC1(input [1:64] in, output [1:56] out);
  assign out[1] = in[57];
  assign out[2] = in[49];
  assign out[3] = in[41];
  assign out[4] = in[33];
  assign out[5] = in[25];
  assign out[6] = in[17];
  assign out[7] = in[9];
  assign out[8] = in[1];
  assign out[9] = in[58];
  assign out[10] = in[50];
  assign out[11] = in[42];
  assign out[12] = in[34];
  assign out[13] = in[26];
  assign out[14] = in[18];
  assign out[15] = in[10];
  assign out[16] = in[2];
  assign out[17] = in[59];
  assign out[18] = in[51];
  assign out[19] = in[43];
  assign out[20] = in[35];
  assign out[21] = in[27];
  assign out[22] = in[19];
  assign out[23] = in[11];
  assign out[24] = in[3];
  assign out[25] = in[60];
  assign out[26] = in[52];
  assign out[27] = in[44];
  assign out[28] = in[36];
  assign out[29] = in[63];
  assign out[30] = in[55];
  assign out[31] = in[47];
  assign out[32] = in[39];
  assign out[33] = in[31];
  assign out[34] = in[23];
  assign out[35] = in[15];
  assign out[36] = in[7];
  assign out[37] = in[62];
  assign out[38] = in[54];
  assign out[39] = in[46];
  assign out[40] = in[38];
  assign out[41] = in[30];
  assign out[42] = in[22];
  assign out[43] = in[14];
  assign out[44] = in[6];
  assign out[45] = in[61];
  assign out[46] = in[53];
  assign out[47] = in[45];
  assign out[48] = in[37];
  assign out[49] = in[29];
  assign out[50] = in[21];
  assign out[51] = in[13];
  assign out[52] = in[5];
  assign out[53] = in[28];
  assign out[54] = in[20];
  assign out[55] = in[12];
  assign out[56] = in[4];
endmodule
module PC2(input [1:56] in, output [1:48] out);
  assign out[1] = in[14];
  assign out[2] = in[17];
  assign out[3] = in[11];
  assign out[4] = in[24];
  assign out[5] = in[1];
  assign out[6] = in[5];
  assign out[7] = in[3];
  assign out[8] = in[28];
  assign out[9] = in[15];
  assign out[10] = in[6];
  assign out[11] = in[21];
  assign out[12] = in[10];
  assign out[13] = in[23];
  assign out[14] = in[19];
  assign out[15] = in[12];
  assign out[16] = in[4];
  assign out[17] = in[26];
  assign out[18] = in[8];
  assign out[19] = in[16];
  assign out[20] = in[7];
  assign out[21] = in[27];
  assign out[22] = in[20];
  assign out[23] = in[13];
  assign out[24] = in[2];
  assign out[25] = in[41];
  assign out[26] = in[52];
  assign out[27] = in[31];
  assign out[28] = in[37];
  assign out[29] = in[47];
  assign out[30] = in[55];
  assign out[31] = in[30];
  assign out[32] = in[40];
  assign out[33] = in[51];
  assign out[34] = in[45];
  assign out[35] = in[33];
  assign out[36] = in[48];
  assign out[37] = in[44];
  assign out[38] = in[49];
  assign out[39] = in[39];
  assign out[40] = in[56];
  assign out[41] = in[34];
  assign out[42] = in[53];
  assign out[43] = in[46];
  assign out[44] = in[42];
  assign out[45] = in[50];
  assign out[46] = in[36];
  assign out[47] = in[29];
  assign out[48] = in[32];
endmodule

module f(input [32:1] R, input [48:1] K, output [32:1] OUT);
  wire [48:1] R_E;
  E E_inst(R, R_E);

  wire [48:1] T = R_E ^ K;

  wire [6:1] S1_in, S2_in, S3_in, S4_in, S5_in, S6_in, S7_in, S8_in;
  assign {S1_in, S2_in, S3_in, S4_in, S5_in, S6_in, S7_in, S8_in} = T;

  wire [4:1] S1_out, S2_out, S3_out, S4_out, S5_out, S6_out, S7_out, S8_out;
  S1 S1_inst(S1_in, S1_out);
  S2 S2_inst(S2_in, S2_out);
  S3 S3_inst(S3_in, S3_out);
  S4 S4_inst(S4_in, S4_out);
  S5 S5_inst(S5_in, S5_out);
  S6 S6_inst(S6_in, S6_out);
  S7 S7_inst(S7_in, S7_out);
  S8 S8_inst(S8_in, S8_out);

  wire [32:1] S_out = {S1_out, S2_out, S3_out, S4_out, S5_out, S6_out, S7_out, S8_out};
  P P_inst(S_out, OUT);
endmodule

module KS_left_shift(input [5:1] level, input [28:1] in, output [28:1] out);
  assign out = (level == 1 || level == 2 || level == 9 || level == 16) ?
                {in[27:1], in[28]} : {in[26:1], in[28:27]};
endmodule

module KS(input [64:1] key, output [48:1] k1,
                            output [48:1] k2,
                            output [48:1] k3,
                            output [48:1] k4,
                            output [48:1] k5,
                            output [48:1] k6,
                            output [48:1] k7,
                            output [48:1] k8,
                            output [48:1] k9,
                            output [48:1] k10,
                            output [48:1] k11,
                            output [48:1] k12,
                            output [48:1] k13,
                            output [48:1] k14,
                            output [48:1] k15,
                            output [48:1] k16);
  wire [56:1] key_pc1;
  PC1 pc1_inst(key, key_pc1);

  wire [28:1] c [0:16];
  wire [28:1] d [0:16];
  wire [48:1] k [1:16];

  assign {c[0], d[0]} = key_pc1;

  genvar i;
  generate
    for (i = 1; i <= 16; i = i + 1) begin : blk
      wire [5:1] j = i;
      KS_left_shift KS_ls_inst1(j, c[i - 1], c[i]);
      KS_left_shift KS_ls_inst2(j, d[i - 1], d[i]);
      PC2 pc2_inst({c[i], d[i]}, k[i]);
    end
  endgenerate

  assign k1 = k[1];
  assign k2 = k[2];
  assign k3 = k[3];
  assign k4 = k[4];
  assign k5 = k[5];
  assign k6 = k[6];
  assign k7 = k[7];
  assign k8 = k[8];
  assign k9 = k[9];
  assign k10 = k[10];
  assign k11 = k[11];
  assign k12 = k[12];
  assign k13 = k[13];
  assign k14 = k[14];
  assign k15 = k[15];
  assign k16 = k[16];
endmodule

module DES_enc(input [64:1] in, input [64:1] key, output [64:1] out);
  wire [64:1] in_ip;
  IP ip_inst(in, in_ip);

  wire [32:1] l [0:16];
  wire [32:1] r [0:16];
  wire [32:1] f_val [1:16];
  assign {l[0], r[0]} = in_ip;

  wire [48:1] k [1:16];
  KS ks_inst(key, k[1], k[2], k[3], k[4], k[5], k[6], k[7], k[8], k[9],
                  k[10], k[11], k[12], k[13], k[14], k[15], k[16]);

  genvar i;
  generate
    for (i = 1; i <= 16; i = i + 1) begin : blk
      assign l[i] = r[i - 1];
      f f_inst(r[i - 1], k[i], f_val[i]);
      assign r[i] = l[i - 1] ^ f_val[i];
    end
  endgenerate

  IP_inv ip_inv_inst({r[16], l[16]}, out);
endmodule

module DES_dec(input [64:1] in, input [64:1] key, output [64:1] out);
  wire [64:1] in_ip;
  IP ip_inst(in, in_ip);

  wire [32:1] l [0:16];
  wire [32:1] r [0:16];
  wire [32:1] f_val [1:16];
  assign {l[0], r[0]} = in_ip;

  wire [48:1] k [1:16];
  KS ks_inst(key, k[16], k[15], k[14], k[13], k[12], k[11], k[10], k[9],
                  k[8], k[7], k[6], k[5], k[4], k[3], k[2], k[1]); // Reverse order

  genvar i;
  generate
    for (i = 1; i <= 16; i = i + 1) begin : blk
      assign l[i] = r[i - 1];
      f f_inst(r[i - 1], k[i], f_val[i]);
      assign r[i] = l[i - 1] ^ f_val[i];
    end
  endgenerate

  IP_inv ip_inv_inst({r[16], l[16]}, out);
endmodule

